module mux4x1 (
   input [3:0] f1;
   input [3:0] f2;
   input [3:0] f3;
   input [3:0] f4;
);
