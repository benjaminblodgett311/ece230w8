module mux4x1 (
    input wire [3:0] sw, 
    output wire led0     
);
  